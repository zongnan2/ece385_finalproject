
module sram_pll (
	clk_clk,
	reset_reset_n,
	sram_clk_clk);	

	input		clk_clk;
	input		reset_reset_n;
	output		sram_clk_clk;
endmodule
